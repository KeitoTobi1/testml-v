module testml

// TODO:Support YAML.
import json

pub type Object =  Null | Integer | Regex | String | Float | Json | Yaml |